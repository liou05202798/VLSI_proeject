* File: freqdiv4_2.pex.netlist
* Created: Mon Jan 13 15:47:11 2020
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "freqdiv4_2.pex.netlist.pex"
.subckt Clock_Divider  CLK_OUT VDD VSS CON1 CON2 CON3 CLK
* 
* CLK	CLK
* CON3	CON3
* CON2	CON2
* CON1	CON1
* VSS	VSS
* VDD	VDD
* CLK_OUT	CLK_OUT
mXI24.MN_inv N_CLK3_XI24.MN_inv_d N_CLK_XI24.MN_inv_g N_VSS_XI24.MN_inv_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=1.07e-12 AS=9.8e-13 PD=3.07e-06
+ PS=2.98e-06
mXI258.MN_inv N_VDD_BAR_XI258.MN_inv_d N_VDD_XI258.MN_inv_g N_VSS_XI258.MN_inv_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI17.X11.MM3 N_DIV7_XI17.X11.MM3_d N_CON1_XI17.X11.MM3_g
+ N_XI17.X11.NET11_XI17.X11.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.225e-13 AS=1.4875e-13 PD=1.79e-06 PS=5.95e-07
mXI17.X11.MM2 N_XI17.X11.NET11_XI17.X11.MM2_d N_CON2_XI17.X11.MM2_g
+ N_XI17.X11.NET7_XI17.X11.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X11.MN_nand3 N_XI17.X11.NET7_XI17.X11.MN_nand3_d
+ N_CON3_XI17.X11.MN_nand3_g N_VSS_XI17.X11.MN_nand3_s N_VSS_XI214.MN_inv_b N_18
+ L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X10.MM3 N_DIV6_XI17.X10.MM3_d N_CON1_XI17.X10.MM3_g
+ N_XI17.X10.NET11_XI17.X10.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.475e-13 AS=1.4875e-13 PD=1.89e-06 PS=5.95e-07
mXI17.X10.MM2 N_XI17.X10.NET11_XI17.X10.MM2_d N_CON2_XI17.X10.MM2_g
+ N_XI17.X10.NET7_XI17.X10.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X10.MN_nand3 N_XI17.X10.NET7_XI17.X10.MN_nand3_d
+ N_XI17.CON3_BAR_XI17.X10.MN_nand3_g N_VSS_XI17.X10.MN_nand3_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X9.MM3 N_DIV5_XI17.X9.MM3_d N_CON1_XI17.X9.MM3_g
+ N_XI17.X9.NET11_XI17.X9.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.2e-13 AS=1.4875e-13 PD=1.78e-06 PS=5.95e-07
mXI17.X9.MM2 N_XI17.X9.NET11_XI17.X9.MM2_d N_XI17.CON2_BAR_XI17.X9.MM2_g
+ N_XI17.X9.NET7_XI17.X9.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X9.MN_nand3 N_XI17.X9.NET7_XI17.X9.MN_nand3_d N_CON3_XI17.X9.MN_nand3_g
+ N_VSS_XI17.X9.MN_nand3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.6e-13 AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X8.MM3 N_DIV4_XI17.X8.MM3_d N_CON1_XI17.X8.MM3_g
+ N_XI17.X8.NET11_XI17.X8.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.375e-13 AS=1.4875e-13 PD=1.85e-06 PS=5.95e-07
mXI17.X8.MM2 N_XI17.X8.NET11_XI17.X8.MM2_d N_XI17.CON2_BAR_XI17.X8.MM2_g
+ N_XI17.X8.NET7_XI17.X8.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X8.MN_nand3 N_XI17.X8.NET7_XI17.X8.MN_nand3_d
+ N_XI17.CON3_BAR_XI17.X8.MN_nand3_g N_VSS_XI17.X8.MN_nand3_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X7.MM3 N_DIV3_XI17.X7.MM3_d N_XI17.CON1_BAR_XI17.X7.MM3_g
+ N_XI17.X7.NET11_XI17.X7.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.225e-13 AS=1.4875e-13 PD=1.79e-06 PS=5.95e-07
mXI17.X7.MM2 N_XI17.X7.NET11_XI17.X7.MM2_d N_CON2_XI17.X7.MM2_g
+ N_XI17.X7.NET7_XI17.X7.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X7.MN_nand3 N_XI17.X7.NET7_XI17.X7.MN_nand3_d N_CON3_XI17.X7.MN_nand3_g
+ N_VSS_XI17.X7.MN_nand3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.6e-13 AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X6.MM3 N_DIV2_XI17.X6.MM3_d N_XI17.CON1_BAR_XI17.X6.MM3_g
+ N_XI17.X6.NET11_XI17.X6.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.175e-13 AS=1.4875e-13 PD=1.77e-06 PS=5.95e-07
mXI17.X6.MM2 N_XI17.X6.NET11_XI17.X6.MM2_d N_CON2_XI17.X6.MM2_g
+ N_XI17.X6.NET7_XI17.X6.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X6.MN_nand3 N_XI17.X6.NET7_XI17.X6.MN_nand3_d
+ N_XI17.CON3_BAR_XI17.X6.MN_nand3_g N_VSS_XI17.X6.MN_nand3_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X5.MM3 N_DIV1_XI17.X5.MM3_d N_XI17.CON1_BAR_XI17.X5.MM3_g
+ N_XI17.X5.NET11_XI17.X5.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.2e-13 AS=1.5875e-13 PD=1.78e-06 PS=6.35e-07
mXI17.X5.MM2 N_XI17.X5.NET11_XI17.X5.MM2_d N_XI17.CON2_BAR_XI17.X5.MM2_g
+ N_XI17.X5.NET7_XI17.X5.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.5875e-13 AS=1.5e-13 PD=6.35e-07 PS=6e-07
mXI17.X5.MN_nand3 N_XI17.X5.NET7_XI17.X5.MN_nand3_d N_CON3_XI17.X5.MN_nand3_g
+ N_VSS_XI17.X5.MN_nand3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.5e-13 AS=2.45e-13 PD=6e-07 PS=1.48e-06
mXI17.X4.MM3 N_XX_XI17.X4.MM3_d N_XI17.CON1_BAR_XI17.X4.MM3_g
+ N_XI17.X4.NET11_XI17.X4.MM3_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=3.15e-13 AS=1.4875e-13 PD=1.76e-06 PS=5.95e-07
mXI17.X4.MM2 N_XI17.X4.NET11_XI17.X4.MM2_d N_XI17.CON2_BAR_XI17.X4.MM2_g
+ N_XI17.X4.NET7_XI17.X4.MM2_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07
+ AD=1.4875e-13 AS=1.6e-13 PD=5.95e-07 PS=6.4e-07
mXI17.X4.MN_nand3 N_XI17.X4.NET7_XI17.X4.MN_nand3_d
+ N_XI17.CON3_BAR_XI17.X4.MN_nand3_g N_VSS_XI17.X4.MN_nand3_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X3.MN_inv N_XI17.CON1_BAR_XI17.X3.MN_inv_d N_CON1_XI17.X3.MN_inv_g
+ N_VSS_XI17.X3.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17.X2.MN_inv N_XI17.CON2_BAR_XI17.X2.MN_inv_d N_CON2_XI17.X2.MN_inv_g
+ N_VSS_XI17.X2.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17.X1.MN_inv N_XI17.CON3_BAR_XI17.X1.MN_inv_d N_CON3_XI17.X1.MN_inv_g
+ N_VSS_XI17.X1.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI24.MP_inv N_CLK3_XI24.MP_inv_d N_CLK_XI24.MP_inv_g N_VDD_XI24.MP_inv_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=6e-06 AD=3.36e-12 AS=2.94e-12
+ PD=7.12e-06 PS=6.98e-06
mXI258.MP_inv N_VDD_BAR_XI258.MP_inv_d N_VDD_XI258.MP_inv_g N_VDD_XI258.MP_inv_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI17.X11.MM5 N_DIV7_XI17.X11.MM5_d N_CON1_XI17.X11.MM5_g N_VDD_XI17.X11.MM5_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.225e-13 AS=1.4875e-13
+ PD=1.79e-06 PS=5.95e-07
mXI17.X11.MM0 N_DIV7_XI17.X11.MM0_d N_CON2_XI17.X11.MM0_g N_VDD_XI17.X11.MM0_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=1.4875e-13
+ PD=6.4e-07 PS=5.95e-07
mXI17.X11.MM4 N_DIV7_XI17.X11.MM4_d N_CON3_XI17.X11.MM4_g N_VDD_XI17.X11.MM4_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X10.MM5 N_DIV6_XI17.X10.MM5_d N_CON1_XI17.X10.MM5_g N_VDD_XI17.X10.MM5_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.475e-13 AS=1.4875e-13
+ PD=1.89e-06 PS=5.95e-07
mXI17.X10.MM0 N_DIV6_XI17.X10.MM0_d N_CON2_XI17.X10.MM0_g N_VDD_XI17.X10.MM0_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=1.4875e-13
+ PD=6.4e-07 PS=5.95e-07
mXI17.X10.MM4 N_DIV6_XI17.X10.MM4_d N_XI17.CON3_BAR_XI17.X10.MM4_g
+ N_VDD_XI17.X10.MM4_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X9.MM5 N_DIV5_XI17.X9.MM5_d N_CON1_XI17.X9.MM5_g N_VDD_XI17.X9.MM5_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.2e-13 AS=1.4875e-13
+ PD=1.78e-06 PS=5.95e-07
mXI17.X9.MM0 N_DIV5_XI17.X9.MM0_d N_XI17.CON2_BAR_XI17.X9.MM0_g
+ N_VDD_XI17.X9.MM0_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=1.4875e-13 PD=6.4e-07 PS=5.95e-07
mXI17.X9.MM4 N_DIV5_XI17.X9.MM4_d N_CON3_XI17.X9.MM4_g N_VDD_XI17.X9.MM4_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X8.MM5 N_DIV4_XI17.X8.MM5_d N_CON1_XI17.X8.MM5_g N_VDD_XI17.X8.MM5_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.375e-13 AS=1.4875e-13
+ PD=1.85e-06 PS=5.95e-07
mXI17.X8.MM0 N_DIV4_XI17.X8.MM0_d N_XI17.CON2_BAR_XI17.X8.MM0_g
+ N_VDD_XI17.X8.MM0_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=1.4875e-13 PD=6.4e-07 PS=5.95e-07
mXI17.X8.MM4 N_DIV4_XI17.X8.MM4_d N_XI17.CON3_BAR_XI17.X8.MM4_g
+ N_VDD_XI17.X8.MM4_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X7.MM5 N_DIV3_XI17.X7.MM5_d N_XI17.CON1_BAR_XI17.X7.MM5_g
+ N_VDD_XI17.X7.MM5_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.225e-13
+ AS=1.4875e-13 PD=1.79e-06 PS=5.95e-07
mXI17.X7.MM0 N_DIV3_XI17.X7.MM0_d N_CON2_XI17.X7.MM0_g N_VDD_XI17.X7.MM0_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=1.4875e-13
+ PD=6.4e-07 PS=5.95e-07
mXI17.X7.MM4 N_DIV3_XI17.X7.MM4_d N_CON3_XI17.X7.MM4_g N_VDD_XI17.X7.MM4_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=2.45e-13 PD=6.4e-07
+ PS=1.48e-06
mXI17.X6.MM5 N_DIV2_XI17.X6.MM5_d N_XI17.CON1_BAR_XI17.X6.MM5_g
+ N_VDD_XI17.X6.MM5_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.175e-13
+ AS=1.4875e-13 PD=1.77e-06 PS=5.95e-07
mXI17.X6.MM0 N_DIV2_XI17.X6.MM0_d N_CON2_XI17.X6.MM0_g N_VDD_XI17.X6.MM0_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13 AS=1.4875e-13
+ PD=6.4e-07 PS=5.95e-07
mXI17.X6.MM4 N_DIV2_XI17.X6.MM4_d N_XI17.CON3_BAR_XI17.X6.MM4_g
+ N_VDD_XI17.X6.MM4_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X5.MM5 N_DIV1_XI17.X5.MM5_d N_XI17.CON1_BAR_XI17.X5.MM5_g
+ N_VDD_XI17.X5.MM5_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.2e-13
+ AS=1.5875e-13 PD=1.78e-06 PS=6.35e-07
mXI17.X5.MM0 N_DIV1_XI17.X5.MM0_d N_XI17.CON2_BAR_XI17.X5.MM0_g
+ N_VDD_XI17.X5.MM0_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.5e-13
+ AS=1.5875e-13 PD=6e-07 PS=6.35e-07
mXI17.X5.MM4 N_DIV1_XI17.X5.MM4_d N_CON3_XI17.X5.MM4_g N_VDD_XI17.X5.MM4_s
+ N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.5e-13 AS=2.45e-13 PD=6e-07
+ PS=1.48e-06
mXI17.X4.MM5 N_XX_XI17.X4.MM5_d N_XI17.CON1_BAR_XI17.X4.MM5_g
+ N_VDD_XI17.X4.MM5_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=3.15e-13
+ AS=1.4875e-13 PD=1.76e-06 PS=5.95e-07
mXI17.X4.MM0 N_XX_XI17.X4.MM0_d N_XI17.CON2_BAR_XI17.X4.MM0_g
+ N_VDD_XI17.X4.MM0_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=1.4875e-13 PD=6.4e-07 PS=5.95e-07
mXI17.X4.MM4 N_XX_XI17.X4.MM4_d N_XI17.CON3_BAR_XI17.X4.MM4_g
+ N_VDD_XI17.X4.MM4_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=1.6e-13
+ AS=2.45e-13 PD=6.4e-07 PS=1.48e-06
mXI17.X3.MP_inv N_XI17.CON1_BAR_XI17.X3.MP_inv_d N_CON1_XI17.X3.MP_inv_g
+ N_VDD_XI17.X3.MP_inv_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17.X2.MP_inv N_XI17.CON2_BAR_XI17.X2.MP_inv_d N_CON2_XI17.X2.MP_inv_g
+ N_VDD_XI17.X2.MP_inv_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17.X1.MP_inv N_XI17.CON3_BAR_XI17.X1.MP_inv_d N_CON3_XI17.X1.MP_inv_g
+ N_VDD_XI17.X1.MP_inv_s N_VDD_XI17.X11.MM5_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI214.MN_inv N_CLK_BY_1_BAR3_XI214.MN_inv_d N_CLK_BY_1_BAR2_XI214.MN_inv_g
+ N_VSS_XI214.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI6.MM0 N_CLK_BY_1_BAR3_XI6.MM0_d N_XI6.NET8_XI6.MM0_g N_CLK_OUT_XI6.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI6.XI0.MN_inv N_XI6.NET8_XI6.XI0.MN_inv_d N_DIV1_XI6.XI0.MN_inv_g
+ N_VSS_XI6.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI214.MP_inv N_CLK_BY_1_BAR3_XI214.MP_inv_d N_CLK_BY_1_BAR2_XI214.MP_inv_g
+ N_VDD_XI214.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI6.MM1 N_CLK_BY_1_BAR3_XI6.MM1_d N_DIV1_XI6.MM1_g N_CLK_OUT_XI6.MM1_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI6.XI0.MP_inv N_XI6.NET8_XI6.XI0.MP_inv_d N_DIV1_XI6.XI0.MP_inv_g
+ N_VDD_XI6.XI0.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI282.MN_inv N_CLK_BY_4_BAR2_XI282.MN_inv_d N_CLK_BY_4_XI282.MN_inv_g
+ N_VSS_XI282.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI13.MM0 N_CLK_BY_4_BAR2_XI13.MM0_d N_XI13.NET8_XI13.MM0_g N_CLK_OUT_XI13.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI13.XI0.MN_inv N_XI13.NET8_XI13.XI0.MN_inv_d N_DIV4_XI13.XI0.MN_inv_g
+ N_VSS_XI13.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI282.MP_inv N_CLK_BY_4_BAR2_XI282.MP_inv_d N_CLK_BY_4_XI282.MP_inv_g
+ N_VDD_XI282.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI13.MM1 N_CLK_BY_4_BAR2_XI13.MM1_d N_DIV4_XI13.MM1_g N_CLK_OUT_XI13.MM1_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI13.XI0.MP_inv N_XI13.NET8_XI13.XI0.MP_inv_d N_DIV4_XI13.XI0.MP_inv_g
+ N_VDD_XI13.XI0.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI278.MN_inv N_CLK_BY_2_BAR3_XI278.MN_inv_d N_CLK_BY_2_BAR2_XI278.MN_inv_g
+ N_VSS_XI278.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI7.MM0 N_CLK_BY_2_BAR3_XI7.MM0_d N_XI7.NET8_XI7.MM0_g N_CLK_OUT_XI7.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI7.XI0.MN_inv N_XI7.NET8_XI7.XI0.MN_inv_d N_DIV2_XI7.XI0.MN_inv_g
+ N_VSS_XI7.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI278.MP_inv N_CLK_BY_2_BAR3_XI278.MP_inv_d N_CLK_BY_2_BAR2_XI278.MP_inv_g
+ N_VDD_XI278.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI7.MM1 N_CLK_BY_2_BAR3_XI7.MM1_d N_DIV2_XI7.MM1_g N_CLK_OUT_XI7.MM1_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI7.XI0.MP_inv N_XI7.NET8_XI7.XI0.MP_inv_d N_DIV2_XI7.XI0.MP_inv_g
+ N_VDD_XI7.XI0.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI262.MN_inv N_CLK_BY_6_BAR2_XI262.MN_inv_d N_CLK_BY_6_XI262.MN_inv_g
+ N_VSS_XI262.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI15.MM0 N_CLK_BY_6_BAR2_XI15.MM0_d N_XI15.NET8_XI15.MM0_g N_CLK_OUT_XI15.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI15.XI0.MN_inv N_XI15.NET8_XI15.XI0.MN_inv_d N_DIV6_XI15.XI0.MN_inv_g
+ N_VSS_XI15.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI262.MP_inv N_CLK_BY_6_BAR2_XI262.MP_inv_d N_CLK_BY_6_XI262.MP_inv_g
+ N_VDD_XI262.MP_inv_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI15.MM1 N_CLK_BY_6_BAR2_XI15.MM1_d N_DIV6_XI15.MM1_g N_CLK_OUT_XI15.MM1_s
+ N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI15.XI0.MP_inv N_XI15.NET8_XI15.XI0.MP_inv_d N_DIV6_XI15.XI0.MP_inv_g
+ N_VDD_XI15.XI0.MP_inv_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI272.MN_inv N_CLK_BY_5_BAR2_XI272.MN_inv_d N_CLK_BY_5_XI272.MN_inv_g
+ N_VSS_XI272.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI14.MM0 N_CLK_BY_5_BAR2_XI14.MM0_d N_XI14.NET8_XI14.MM0_g N_CLK_OUT_XI14.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI14.XI0.MN_inv N_XI14.NET8_XI14.XI0.MN_inv_d N_DIV5_XI14.XI0.MN_inv_g
+ N_VSS_XI14.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI272.MP_inv N_CLK_BY_5_BAR2_XI272.MP_inv_d N_CLK_BY_5_XI272.MP_inv_g
+ N_VDD_XI272.MP_inv_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI14.MM1 N_CLK_BY_5_BAR2_XI14.MM1_d N_DIV5_XI14.MM1_g N_CLK_OUT_XI14.MM1_s
+ N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI14.XI0.MP_inv N_XI14.NET8_XI14.XI0.MP_inv_d N_DIV5_XI14.XI0.MP_inv_g
+ N_VDD_XI14.XI0.MP_inv_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI254.MN_inv N_VDD_BAR2_XI254.MN_inv_d N_VDD_BAR_XI254.MN_inv_g
+ N_VSS_XI254.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI5.MM0 N_VDD_BAR2_XI5.MM0_d N_XI5.NET8_XI5.MM0_g N_CLK_OUT_XI5.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI5.XI0.MN_inv N_XI5.NET8_XI5.XI0.MN_inv_d N_XX_XI5.XI0.MN_inv_g
+ N_VSS_XI5.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI254.MP_inv N_VDD_BAR2_XI254.MP_inv_d N_VDD_BAR_XI254.MP_inv_g
+ N_VDD_XI254.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI5.MM1 N_VDD_BAR2_XI5.MM1_d N_XX_XI5.MM1_g N_CLK_OUT_XI5.MM1_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI5.XI0.MP_inv N_XI5.NET8_XI5.XI0.MP_inv_d N_XX_XI5.XI0.MP_inv_g
+ N_VDD_XI5.XI0.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI298.MN_inv N_CLK_BY_3_BAR3_XI298.MN_inv_d N_CLK_BY_3_BAR2_XI298.MN_inv_g
+ N_VSS_XI298.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI8.MM0 N_CLK_BY_3_BAR3_XI8.MM0_d N_XI8.NET8_XI8.MM0_g N_CLK_OUT_XI8.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI8.XI0.MN_inv N_XI8.NET8_XI8.XI0.MN_inv_d N_DIV3_XI8.XI0.MN_inv_g
+ N_VSS_XI8.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI298.MP_inv N_CLK_BY_3_BAR3_XI298.MP_inv_d N_CLK_BY_3_BAR2_XI298.MP_inv_g
+ N_VDD_XI298.MP_inv_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI8.MM1 N_CLK_BY_3_BAR3_XI8.MM1_d N_DIV3_XI8.MM1_g N_CLK_OUT_XI8.MM1_s
+ N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI8.XI0.MP_inv N_XI8.NET8_XI8.XI0.MP_inv_d N_DIV3_XI8.XI0.MP_inv_g
+ N_VDD_XI8.XI0.MP_inv_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI252.MN_inv N_CLK_BY_7_BAR2_XI252.MN_inv_d N_CLK_BY_7_XI252.MN_inv_g
+ N_VSS_XI252.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13
+ AS=9.88e-13 PD=5.15e-07 PS=2.988e-06
mXI16.MM0 N_CLK_BY_7_BAR2_XI16.MM0_d N_XI16.NET8_XI16.MM0_g N_CLK_OUT_XI16.MM0_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=5.15e-13 AS=1.012e-12
+ PD=5.15e-07 PS=3.012e-06
mXI16.XI0.MN_inv N_XI16.NET8_XI16.XI0.MN_inv_d N_DIV7_XI16.XI0.MN_inv_g
+ N_VSS_XI16.XI0.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=9.8e-13
+ AS=1.012e-12 PD=2.98e-06 PS=3.012e-06
mXI252.MP_inv N_CLK_BY_7_BAR2_XI252.MP_inv_d N_CLK_BY_7_XI252.MP_inv_g
+ N_VDD_XI252.MP_inv_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12
+ AS=1.976e-12 PD=5.15e-07 PS=4.988e-06
mXI16.MM1 N_CLK_BY_7_BAR2_XI16.MM1_d N_DIV7_XI16.MM1_g N_CLK_OUT_XI16.MM1_s
+ N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=4e-06 AD=1.03e-12 AS=2.016e-12
+ PD=5.15e-07 PS=5.008e-06
mXI16.XI0.MP_inv N_XI16.NET8_XI16.XI0.MP_inv_d N_DIV7_XI16.XI0.MP_inv_g
+ N_VDD_XI16.XI0.MP_inv_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=4e-06
+ AD=1.976e-12 AS=2.016e-12 PD=4.988e-06 PS=5.008e-06
mXI19.XI0.MM8 N_XI19.XI0.NET15_XI19.XI0.MM8_d N_XI19.NET8_XI19.XI0.MM8_g
+ N_VSS_XI19.XI0.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI19.XI0.MM9 N_XI19.XI0.NET11_XI19.XI0.MM9_d N_CLK3_XI19.XI0.MM9_g
+ N_VSS_XI19.XI0.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI19.XI0.MM5 N_XI19.XI0.NET27_XI19.XI0.MM5_d N_XI19.XI0.NET15_XI19.XI0.MM5_g
+ N_XI19.XI0.NET11_XI19.XI0.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI19.XI0.MM10 N_XI19.XI0.NET7_XI19.XI0.MM10_d N_XI19.XI0.NET27_XI19.XI0.MM10_g
+ N_VSS_XI19.XI0.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI19.XI0.MM6 N_XI19.NET25_XI19.XI0.MM6_d N_CLK3_XI19.XI0.MM6_g
+ N_XI19.XI0.NET7_XI19.XI0.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI19.XI0.MM7 N_XI19.NET7_XI19.XI0.MM7_d N_XI19.NET25_XI19.XI0.MM7_g
+ N_VSS_XI19.XI0.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI19.XI0.MM0 N_XI19.XI0.NET34_XI19.XI0.MM0_d N_XI19.NET8_XI19.XI0.MM0_g
+ N_VDD_XI19.XI0.MM0_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI19.XI0.MM4 N_XI19.XI0.NET15_XI19.XI0.MM4_d N_CLK3_XI19.XI0.MM4_g
+ N_XI19.XI0.NET34_XI19.XI0.MM4_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI19.XI0.MM1 N_XI19.XI0.NET27_XI19.XI0.MM1_d N_CLK3_XI19.XI0.MM1_g
+ N_VDD_XI19.XI0.MM1_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI19.XI0.MM2 N_XI19.NET25_XI19.XI0.MM2_d N_XI19.XI0.NET27_XI19.XI0.MM2_g
+ N_VDD_XI19.XI0.MM2_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI19.XI0.MM3 N_XI19.NET7_XI19.XI0.MM3_d N_XI19.NET25_XI19.XI0.MM3_g
+ N_VDD_XI19.XI0.MM3_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI21.XI0.MM8 N_XI21.XI0.NET15_XI21.XI0.MM8_d N_XI21.NET7_XI21.XI0.MM8_g
+ N_VSS_XI21.XI0.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI21.XI0.MM9 N_XI21.XI0.NET11_XI21.XI0.MM9_d N_CLK3_XI21.XI0.MM9_g
+ N_VSS_XI21.XI0.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI21.XI0.MM5 N_XI21.XI0.NET27_XI21.XI0.MM5_d N_XI21.XI0.NET15_XI21.XI0.MM5_g
+ N_XI21.XI0.NET11_XI21.XI0.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI21.XI0.MM10 N_XI21.XI0.NET7_XI21.XI0.MM10_d N_XI21.XI0.NET27_XI21.XI0.MM10_g
+ N_VSS_XI21.XI0.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI21.XI0.MM6 N_XI21.NET30_XI21.XI0.MM6_d N_CLK3_XI21.XI0.MM6_g
+ N_XI21.XI0.NET7_XI21.XI0.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI21.XI0.MM7 N_XI21.NET31_XI21.XI0.MM7_d N_XI21.NET30_XI21.XI0.MM7_g
+ N_VSS_XI21.XI0.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI21.XI0.MM0 N_XI21.XI0.NET34_XI21.XI0.MM0_d N_XI21.NET7_XI21.XI0.MM0_g
+ N_VDD_XI21.XI0.MM0_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI21.XI0.MM4 N_XI21.XI0.NET15_XI21.XI0.MM4_d N_CLK3_XI21.XI0.MM4_g
+ N_XI21.XI0.NET34_XI21.XI0.MM4_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI21.XI0.MM1 N_XI21.XI0.NET27_XI21.XI0.MM1_d N_CLK3_XI21.XI0.MM1_g
+ N_VDD_XI21.XI0.MM1_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI21.XI0.MM2 N_XI21.NET30_XI21.XI0.MM2_d N_XI21.XI0.NET27_XI21.XI0.MM2_g
+ N_VDD_XI21.XI0.MM2_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI21.XI0.MM3 N_XI21.NET31_XI21.XI0.MM3_d N_XI21.NET30_XI21.XI0.MM3_g
+ N_VDD_XI21.XI0.MM3_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI20.XI0.MM8 N_XI20.XI0.NET15_XI20.XI0.MM8_d N_XI20.NET7_XI20.XI0.MM8_g
+ N_VSS_XI20.XI0.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI20.XI0.MM9 N_XI20.XI0.NET11_XI20.XI0.MM9_d N_CLK3_XI20.XI0.MM9_g
+ N_VSS_XI20.XI0.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI20.XI0.MM5 N_XI20.XI0.NET27_XI20.XI0.MM5_d N_XI20.XI0.NET15_XI20.XI0.MM5_g
+ N_XI20.XI0.NET11_XI20.XI0.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI20.XI0.MM10 N_XI20.XI0.NET7_XI20.XI0.MM10_d N_XI20.XI0.NET27_XI20.XI0.MM10_g
+ N_VSS_XI20.XI0.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI20.XI0.MM6 N_XI20.NET24_XI20.XI0.MM6_d N_CLK3_XI20.XI0.MM6_g
+ N_XI20.XI0.NET7_XI20.XI0.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI20.XI0.MM7 N_XI20.NET25_XI20.XI0.MM7_d N_XI20.NET24_XI20.XI0.MM7_g
+ N_VSS_XI20.XI0.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI20.XI0.MM0 N_XI20.XI0.NET34_XI20.XI0.MM0_d N_XI20.NET7_XI20.XI0.MM0_g
+ N_VDD_XI20.XI0.MM0_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI20.XI0.MM4 N_XI20.XI0.NET15_XI20.XI0.MM4_d N_CLK3_XI20.XI0.MM4_g
+ N_XI20.XI0.NET34_XI20.XI0.MM4_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI20.XI0.MM1 N_XI20.XI0.NET27_XI20.XI0.MM1_d N_CLK3_XI20.XI0.MM1_g
+ N_VDD_XI20.XI0.MM1_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI20.XI0.MM2 N_XI20.NET24_XI20.XI0.MM2_d N_XI20.XI0.NET27_XI20.XI0.MM2_g
+ N_VDD_XI20.XI0.MM2_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI20.XI0.MM3 N_XI20.NET25_XI20.XI0.MM3_d N_XI20.NET24_XI20.XI0.MM3_g
+ N_VDD_XI20.XI0.MM3_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI21.XI1.MM8 N_XI21.XI1.NET15_XI21.XI1.MM8_d N_XI21.NET31_XI21.XI1.MM8_g
+ N_VSS_XI21.XI1.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI21.XI1.MM9 N_XI21.XI1.NET11_XI21.XI1.MM9_d N_CLK3_XI21.XI1.MM9_g
+ N_VSS_XI21.XI1.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI21.XI1.MM5 N_XI21.XI1.NET27_XI21.XI1.MM5_d N_XI21.XI1.NET15_XI21.XI1.MM5_g
+ N_XI21.XI1.NET11_XI21.XI1.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI21.XI1.MM10 N_XI21.XI1.NET7_XI21.XI1.MM10_d N_XI21.XI1.NET27_XI21.XI1.MM10_g
+ N_VSS_XI21.XI1.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI21.XI1.MM6 N_XI21.NET24_XI21.XI1.MM6_d N_CLK3_XI21.XI1.MM6_g
+ N_XI21.XI1.NET7_XI21.XI1.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI21.XI1.MM7 N_XI21.NET25_XI21.XI1.MM7_d N_XI21.NET24_XI21.XI1.MM7_g
+ N_VSS_XI21.XI1.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI21.XI1.MM0 N_XI21.XI1.NET34_XI21.XI1.MM0_d N_XI21.NET31_XI21.XI1.MM0_g
+ N_VDD_XI21.XI1.MM0_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI21.XI1.MM4 N_XI21.XI1.NET15_XI21.XI1.MM4_d N_CLK3_XI21.XI1.MM4_g
+ N_XI21.XI1.NET34_XI21.XI1.MM4_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI21.XI1.MM1 N_XI21.XI1.NET27_XI21.XI1.MM1_d N_CLK3_XI21.XI1.MM1_g
+ N_VDD_XI21.XI1.MM1_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI21.XI1.MM2 N_XI21.NET24_XI21.XI1.MM2_d N_XI21.XI1.NET27_XI21.XI1.MM2_g
+ N_VDD_XI21.XI1.MM2_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI21.XI1.MM3 N_XI21.NET25_XI21.XI1.MM3_d N_XI21.NET24_XI21.XI1.MM3_g
+ N_VDD_XI21.XI1.MM3_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI18.XOUT_clk.MM8 N_XI18.XOUT_CLK.NET15_XI18.XOUT_clk.MM8_d
+ N_XI18.NET13_XI18.XOUT_clk.MM8_g N_VSS_XI18.XOUT_clk.MM8_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13 AS=5.05e-13
+ PD=2.07e-06 PS=2.01e-06
mXI18.XOUT_clk.MM9 N_XI18.XOUT_CLK.NET11_XI18.XOUT_clk.MM9_d
+ N_CLK3_XI18.XOUT_clk.MM9_g N_VSS_XI18.XOUT_clk.MM9_s N_VSS_XI214.MN_inv_b N_18
+ L=1.8e-07 W=1e-06 AD=2.075e-13 AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI18.XOUT_clk.MM5 N_XI18.XOUT_CLK.NET27_XI18.XOUT_clk.MM5_d
+ N_XI18.XOUT_CLK.NET15_XI18.XOUT_clk.MM5_g
+ N_XI18.XOUT_CLK.NET11_XI18.XOUT_clk.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07
+ W=1e-06 AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI18.XOUT_clk.MM10 N_XI18.XOUT_CLK.NET7_XI18.XOUT_clk.MM10_d
+ N_XI18.XOUT_CLK.NET27_XI18.XOUT_clk.MM10_g N_VSS_XI18.XOUT_clk.MM10_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13 AS=5.4e-13
+ PD=4.75e-07 PS=2.08e-06
mXI18.XOUT_clk.MM6 N_XI18.NET13_XI18.XOUT_clk.MM6_d N_CLK3_XI18.XOUT_clk.MM6_g
+ N_XI18.XOUT_CLK.NET7_XI18.XOUT_clk.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07
+ W=1e-06 AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI18.XOUT_clk.MM7 N_CLK_BY_2_XI18.XOUT_clk.MM7_d
+ N_XI18.NET13_XI18.XOUT_clk.MM7_g N_VSS_XI18.XOUT_clk.MM7_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13 AS=5.3e-13 PD=2.02e-06
+ PS=2.06e-06
mXI18.XOUT_clk.MM0 N_XI18.XOUT_CLK.NET34_XI18.XOUT_clk.MM0_d
+ N_XI18.NET13_XI18.XOUT_clk.MM0_g N_VDD_XI18.XOUT_clk.MM0_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13 AS=1.03e-12
+ PD=3.25e-07 PS=3.03e-06
mXI18.XOUT_clk.MM4 N_XI18.XOUT_CLK.NET15_XI18.XOUT_clk.MM4_d
+ N_CLK3_XI18.XOUT_clk.MM4_g N_XI18.XOUT_CLK.NET34_XI18.XOUT_clk.MM4_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.83e-12 AS=3.25e-13
+ PD=3.83e-06 PS=3.25e-07
mXI18.XOUT_clk.MM1 N_XI18.XOUT_CLK.NET27_XI18.XOUT_clk.MM1_d
+ N_CLK3_XI18.XOUT_clk.MM1_g N_VDD_XI18.XOUT_clk.MM1_s N_VDD_XI214.MP_inv_b P_18
+ L=1.8e-07 W=2e-06 AD=1.37e-12 AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI18.XOUT_clk.MM2 N_XI18.NET13_XI18.XOUT_clk.MM2_d
+ N_XI18.XOUT_CLK.NET27_XI18.XOUT_clk.MM2_g N_VDD_XI18.XOUT_clk.MM2_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12 AS=1.08e-12 PD=3e-06
+ PS=3.08e-06
mXI18.XOUT_clk.MM3 N_CLK_BY_2_XI18.XOUT_clk.MM3_d
+ N_XI18.NET13_XI18.XOUT_clk.MM3_g N_VDD_XI18.XOUT_clk.MM3_s
+ N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12 AS=1.06e-12
+ PD=3.02e-06 PS=3.06e-06
mXI18.XI0.MM8 N_XI18.XI0.NET15_XI18.XI0.MM8_d N_XI18.NET7_XI18.XI0.MM8_g
+ N_VSS_XI18.XI0.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI18.XI0.MM9 N_XI18.XI0.NET11_XI18.XI0.MM9_d N_XI18.NET13_XI18.XI0.MM9_g
+ N_VSS_XI18.XI0.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI18.XI0.MM5 N_XI18.XI0.NET27_XI18.XI0.MM5_d N_XI18.XI0.NET15_XI18.XI0.MM5_g
+ N_XI18.XI0.NET11_XI18.XI0.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI18.XI0.MM10 N_XI18.XI0.NET7_XI18.XI0.MM10_d N_XI18.XI0.NET27_XI18.XI0.MM10_g
+ N_VSS_XI18.XI0.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI18.XI0.MM6 N_XI18.NET7_XI18.XI0.MM6_d N_XI18.NET13_XI18.XI0.MM6_g
+ N_XI18.XI0.NET7_XI18.XI0.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI18.XI0.MM7 N_CLK_BY_4_XI18.XI0.MM7_d N_XI18.NET7_XI18.XI0.MM7_g
+ N_VSS_XI18.XI0.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI18.XI0.MM0 N_XI18.XI0.NET34_XI18.XI0.MM0_d N_XI18.NET7_XI18.XI0.MM0_g
+ N_VDD_XI18.XI0.MM0_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI18.XI0.MM4 N_XI18.XI0.NET15_XI18.XI0.MM4_d N_XI18.NET13_XI18.XI0.MM4_g
+ N_XI18.XI0.NET34_XI18.XI0.MM4_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI18.XI0.MM1 N_XI18.XI0.NET27_XI18.XI0.MM1_d N_XI18.NET13_XI18.XI0.MM1_g
+ N_VDD_XI18.XI0.MM1_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI18.XI0.MM2 N_XI18.NET7_XI18.XI0.MM2_d N_XI18.XI0.NET27_XI18.XI0.MM2_g
+ N_VDD_XI18.XI0.MM2_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI18.XI0.MM3 N_CLK_BY_4_XI18.XI0.MM3_d N_XI18.NET7_XI18.XI0.MM3_g
+ N_VDD_XI18.XI0.MM3_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI19.XI1.MM8 N_XI19.XI1.NET15_XI19.XI1.MM8_d N_XI19.NET7_XI19.XI1.MM8_g
+ N_VSS_XI19.XI1.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI19.XI1.MM9 N_XI19.XI1.NET11_XI19.XI1.MM9_d N_CLK3_XI19.XI1.MM9_g
+ N_VSS_XI19.XI1.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI19.XI1.MM5 N_XI19.XI1.NET27_XI19.XI1.MM5_d N_XI19.XI1.NET15_XI19.XI1.MM5_g
+ N_XI19.XI1.NET11_XI19.XI1.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI19.XI1.MM10 N_XI19.XI1.NET7_XI19.XI1.MM10_d N_XI19.XI1.NET27_XI19.XI1.MM10_g
+ N_VSS_XI19.XI1.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI19.XI1.MM6 N_XI19.NET19_XI19.XI1.MM6_d N_CLK3_XI19.XI1.MM6_g
+ N_XI19.XI1.NET7_XI19.XI1.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI19.XI1.MM7 N_CLK_BY_3_XI19.XI1.MM7_d N_XI19.NET19_XI19.XI1.MM7_g
+ N_VSS_XI19.XI1.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI19.XI1.MM0 N_XI19.XI1.NET34_XI19.XI1.MM0_d N_XI19.NET7_XI19.XI1.MM0_g
+ N_VDD_XI19.XI1.MM0_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI19.XI1.MM4 N_XI19.XI1.NET15_XI19.XI1.MM4_d N_CLK3_XI19.XI1.MM4_g
+ N_XI19.XI1.NET34_XI19.XI1.MM4_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI19.XI1.MM1 N_XI19.XI1.NET27_XI19.XI1.MM1_d N_CLK3_XI19.XI1.MM1_g
+ N_VDD_XI19.XI1.MM1_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI19.XI1.MM2 N_XI19.NET19_XI19.XI1.MM2_d N_XI19.XI1.NET27_XI19.XI1.MM2_g
+ N_VDD_XI19.XI1.MM2_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI19.XI1.MM3 N_CLK_BY_3_XI19.XI1.MM3_d N_XI19.NET19_XI19.XI1.MM3_g
+ N_VDD_XI19.XI1.MM3_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI19.XI2.MM8 N_XI19.XI2.NET15_XI19.XI2.MM8_d N_XI19.NET034_XI19.XI2.MM8_g
+ N_VSS_XI19.XI2.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI19.XI2.MM9 N_XI19.XI2.NET11_XI19.XI2.MM9_d N_CLK_BY_3_XI19.XI2.MM9_g
+ N_VSS_XI19.XI2.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI19.XI2.MM5 N_XI19.XI2.NET27_XI19.XI2.MM5_d N_XI19.XI2.NET15_XI19.XI2.MM5_g
+ N_XI19.XI2.NET11_XI19.XI2.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI19.XI2.MM10 N_XI19.XI2.NET7_XI19.XI2.MM10_d N_XI19.XI2.NET27_XI19.XI2.MM10_g
+ N_VSS_XI19.XI2.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI19.XI2.MM6 N_XI19.NET034_XI19.XI2.MM6_d N_CLK_BY_3_XI19.XI2.MM6_g
+ N_XI19.XI2.NET7_XI19.XI2.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI19.XI2.MM7 N_CLK_BY_6_XI19.XI2.MM7_d N_XI19.NET034_XI19.XI2.MM7_g
+ N_VSS_XI19.XI2.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI19.XI2.MM0 N_XI19.XI2.NET34_XI19.XI2.MM0_d N_XI19.NET034_XI19.XI2.MM0_g
+ N_VDD_XI19.XI2.MM0_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI19.XI2.MM4 N_XI19.XI2.NET15_XI19.XI2.MM4_d N_CLK_BY_3_XI19.XI2.MM4_g
+ N_XI19.XI2.NET34_XI19.XI2.MM4_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI19.XI2.MM1 N_XI19.XI2.NET27_XI19.XI2.MM1_d N_CLK_BY_3_XI19.XI2.MM1_g
+ N_VDD_XI19.XI2.MM1_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI19.XI2.MM2 N_XI19.NET034_XI19.XI2.MM2_d N_XI19.XI2.NET27_XI19.XI2.MM2_g
+ N_VDD_XI19.XI2.MM2_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI19.XI2.MM3 N_CLK_BY_6_XI19.XI2.MM3_d N_XI19.NET034_XI19.XI2.MM3_g
+ N_VDD_XI19.XI2.MM3_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI20.XI1.MM8 N_XI20.XI1.NET15_XI20.XI1.MM8_d N_XI20.NET25_XI20.XI1.MM8_g
+ N_VSS_XI20.XI1.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI20.XI1.MM9 N_XI20.XI1.NET11_XI20.XI1.MM9_d N_CLK3_XI20.XI1.MM9_g
+ N_VSS_XI20.XI1.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI20.XI1.MM5 N_XI20.XI1.NET27_XI20.XI1.MM5_d N_XI20.XI1.NET15_XI20.XI1.MM5_g
+ N_XI20.XI1.NET11_XI20.XI1.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI20.XI1.MM10 N_XI20.XI1.NET7_XI20.XI1.MM10_d N_XI20.XI1.NET27_XI20.XI1.MM10_g
+ N_VSS_XI20.XI1.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI20.XI1.MM6 N_XI20.NET18_XI20.XI1.MM6_d N_CLK3_XI20.XI1.MM6_g
+ N_XI20.XI1.NET7_XI20.XI1.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI20.XI1.MM7 N_XI20.NET6_XI20.XI1.MM7_d N_XI20.NET18_XI20.XI1.MM7_g
+ N_VSS_XI20.XI1.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI20.XI1.MM0 N_XI20.XI1.NET34_XI20.XI1.MM0_d N_XI20.NET25_XI20.XI1.MM0_g
+ N_VDD_XI20.XI1.MM0_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI20.XI1.MM4 N_XI20.XI1.NET15_XI20.XI1.MM4_d N_CLK3_XI20.XI1.MM4_g
+ N_XI20.XI1.NET34_XI20.XI1.MM4_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI20.XI1.MM1 N_XI20.XI1.NET27_XI20.XI1.MM1_d N_CLK3_XI20.XI1.MM1_g
+ N_VDD_XI20.XI1.MM1_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI20.XI1.MM2 N_XI20.NET18_XI20.XI1.MM2_d N_XI20.XI1.NET27_XI20.XI1.MM2_g
+ N_VDD_XI20.XI1.MM2_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI20.XI1.MM3 N_XI20.NET6_XI20.XI1.MM3_d N_XI20.NET18_XI20.XI1.MM3_g
+ N_VDD_XI20.XI1.MM3_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI20.XI2.MM8 N_XI20.XI2.NET15_XI20.XI2.MM8_d N_XI20.NET6_XI20.XI2.MM8_g
+ N_VSS_XI20.XI2.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI20.XI2.MM9 N_XI20.XI2.NET11_XI20.XI2.MM9_d N_CLK3_XI20.XI2.MM9_g
+ N_VSS_XI20.XI2.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI20.XI2.MM5 N_XI20.XI2.NET27_XI20.XI2.MM5_d N_XI20.XI2.NET15_XI20.XI2.MM5_g
+ N_XI20.XI2.NET11_XI20.XI2.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI20.XI2.MM10 N_XI20.XI2.NET7_XI20.XI2.MM10_d N_XI20.XI2.NET27_XI20.XI2.MM10_g
+ N_VSS_XI20.XI2.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI20.XI2.MM6 N_XI20.NET12_XI20.XI2.MM6_d N_CLK3_XI20.XI2.MM6_g
+ N_XI20.XI2.NET7_XI20.XI2.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI20.XI2.MM7 N_CLK_BY_5_XI20.XI2.MM7_d N_XI20.NET12_XI20.XI2.MM7_g
+ N_VSS_XI20.XI2.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI20.XI2.MM0 N_XI20.XI2.NET34_XI20.XI2.MM0_d N_XI20.NET6_XI20.XI2.MM0_g
+ N_VDD_XI20.XI2.MM0_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI20.XI2.MM4 N_XI20.XI2.NET15_XI20.XI2.MM4_d N_CLK3_XI20.XI2.MM4_g
+ N_XI20.XI2.NET34_XI20.XI2.MM4_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI20.XI2.MM1 N_XI20.XI2.NET27_XI20.XI2.MM1_d N_CLK3_XI20.XI2.MM1_g
+ N_VDD_XI20.XI2.MM1_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI20.XI2.MM2 N_XI20.NET12_XI20.XI2.MM2_d N_XI20.XI2.NET27_XI20.XI2.MM2_g
+ N_VDD_XI20.XI2.MM2_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI20.XI2.MM3 N_CLK_BY_5_XI20.XI2.MM3_d N_XI20.NET12_XI20.XI2.MM3_g
+ N_VDD_XI20.XI2.MM3_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI21.XI2.MM8 N_XI21.XI2.NET15_XI21.XI2.MM8_d N_XI21.NET25_XI21.XI2.MM8_g
+ N_VSS_XI21.XI2.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI21.XI2.MM9 N_XI21.XI2.NET11_XI21.XI2.MM9_d N_CLK3_XI21.XI2.MM9_g
+ N_VSS_XI21.XI2.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI21.XI2.MM5 N_XI21.XI2.NET27_XI21.XI2.MM5_d N_XI21.XI2.NET15_XI21.XI2.MM5_g
+ N_XI21.XI2.NET11_XI21.XI2.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI21.XI2.MM10 N_XI21.XI2.NET7_XI21.XI2.MM10_d N_XI21.XI2.NET27_XI21.XI2.MM10_g
+ N_VSS_XI21.XI2.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI21.XI2.MM6 N_XI21.NET18_XI21.XI2.MM6_d N_CLK3_XI21.XI2.MM6_g
+ N_XI21.XI2.NET7_XI21.XI2.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI21.XI2.MM7 N_XI21.NET6_XI21.XI2.MM7_d N_XI21.NET18_XI21.XI2.MM7_g
+ N_VSS_XI21.XI2.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI21.XI2.MM0 N_XI21.XI2.NET34_XI21.XI2.MM0_d N_XI21.NET25_XI21.XI2.MM0_g
+ N_VDD_XI21.XI2.MM0_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI21.XI2.MM4 N_XI21.XI2.NET15_XI21.XI2.MM4_d N_CLK3_XI21.XI2.MM4_g
+ N_XI21.XI2.NET34_XI21.XI2.MM4_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI21.XI2.MM1 N_XI21.XI2.NET27_XI21.XI2.MM1_d N_CLK3_XI21.XI2.MM1_g
+ N_VDD_XI21.XI2.MM1_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI21.XI2.MM2 N_XI21.NET18_XI21.XI2.MM2_d N_XI21.XI2.NET27_XI21.XI2.MM2_g
+ N_VDD_XI21.XI2.MM2_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI21.XI2.MM3 N_XI21.NET6_XI21.XI2.MM3_d N_XI21.NET18_XI21.XI2.MM3_g
+ N_VDD_XI21.XI2.MM3_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI21.XI3.MM8 N_XI21.XI3.NET15_XI21.XI3.MM8_d N_XI21.NET6_XI21.XI3.MM8_g
+ N_VSS_XI21.XI3.MM8_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.35e-13
+ AS=5.05e-13 PD=2.07e-06 PS=2.01e-06
mXI21.XI3.MM9 N_XI21.XI3.NET11_XI21.XI3.MM9_d N_CLK3_XI21.XI3.MM9_g
+ N_VSS_XI21.XI3.MM9_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.075e-13
+ AS=6e-13 PD=4.15e-07 PS=2.2e-06
mXI21.XI3.MM5 N_XI21.XI3.NET27_XI21.XI3.MM5_d N_XI21.XI3.NET15_XI21.XI3.MM5_g
+ N_XI21.XI3.NET11_XI21.XI3.MM5_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=8.6e-13 AS=2.075e-13 PD=2.72e-06 PS=4.15e-07
mXI21.XI3.MM10 N_XI21.XI3.NET7_XI21.XI3.MM10_d N_XI21.XI3.NET27_XI21.XI3.MM10_g
+ N_VSS_XI21.XI3.MM10_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=2.375e-13
+ AS=5.4e-13 PD=4.75e-07 PS=2.08e-06
mXI21.XI3.MM6 N_XI21.NET12_XI21.XI3.MM6_d N_CLK3_XI21.XI3.MM6_g
+ N_XI21.XI3.NET7_XI21.XI3.MM6_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06
+ AD=7.55e-13 AS=2.375e-13 PD=2.51e-06 PS=4.75e-07
mXI21.XI3.MM7 N_CLK_BY_7_XI21.XI3.MM7_d N_XI21.NET12_XI21.XI3.MM7_g
+ N_VSS_XI21.XI3.MM7_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=1e-06 AD=5.1e-13
+ AS=5.3e-13 PD=2.02e-06 PS=2.06e-06
mXI21.XI3.MM0 N_XI21.XI3.NET34_XI21.XI3.MM0_d N_XI21.NET6_XI21.XI3.MM0_g
+ N_VDD_XI21.XI3.MM0_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=3.25e-13
+ AS=1.03e-12 PD=3.25e-07 PS=3.03e-06
mXI21.XI3.MM4 N_XI21.XI3.NET15_XI21.XI3.MM4_d N_CLK3_XI21.XI3.MM4_g
+ N_XI21.XI3.NET34_XI21.XI3.MM4_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=1.83e-12 AS=3.25e-13 PD=3.83e-06 PS=3.25e-07
mXI21.XI3.MM1 N_XI21.XI3.NET27_XI21.XI3.MM1_d N_CLK3_XI21.XI3.MM1_g
+ N_VDD_XI21.XI3.MM1_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.37e-12
+ AS=1.04e-12 PD=3.37e-06 PS=3.04e-06
mXI21.XI3.MM2 N_XI21.NET12_XI21.XI3.MM2_d N_XI21.XI3.NET27_XI21.XI3.MM2_g
+ N_VDD_XI21.XI3.MM2_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1e-12
+ AS=1.08e-12 PD=3e-06 PS=3.08e-06
mXI21.XI3.MM3 N_CLK_BY_7_XI21.XI3.MM3_d N_XI21.NET12_XI21.XI3.MM3_g
+ N_VDD_XI21.XI3.MM3_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=1.02e-12
+ AS=1.06e-12 PD=3.02e-06 PS=3.06e-06
mXI19.Xr.MN_nand2 N_XI19.XR.NET6_XI19.Xr.MN_nand2_d
+ N_XI19.NET7_XI19.Xr.MN_nand2_g N_VSS_XI19.Xr.MN_nand2_s N_VSS_XI214.MN_inv_b
+ N_18 L=1.8e-07 W=2e-06 AD=7.55e-13 AS=1.24e-12 PD=7.55e-07 PS=3.24e-06
mXI19.Xr.MM1 N_XI19.NET8_XI19.Xr.MM1_d N_CLK_BY_3_XI19.Xr.MM1_g
+ N_XI19.XR.NET6_XI19.Xr.MM1_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06
+ AD=1.59e-12 AS=7.55e-13 PD=3.59e-06 PS=7.55e-07
mXI19.Xr.MP_nand2 N_XI19.NET8_XI19.Xr.MP_nand2_d N_XI19.NET7_XI19.Xr.MP_nand2_g
+ N_VDD_XI19.Xr.MP_nand2_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06
+ AD=7.55e-13 AS=1.22e-12 PD=7.55e-07 PS=3.22e-06
mXI19.Xr.MM0 N_XI19.NET8_XI19.Xr.MM0_d N_CLK_BY_3_XI19.Xr.MM0_g
+ N_VDD_XI19.Xr.MM0_s N_VDD_XI262.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=7.55e-13
+ AS=1.38e-12 PD=7.55e-07 PS=3.38e-06
mXI20.XI3.MM1 N_XI20.XI3.NET6_XI20.XI3.MM1_d N_CLK_BY_5_XI20.XI3.MM1_g
+ N_VSS_XI20.XI3.MM1_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=7.55e-13
+ AS=1.24e-12 PD=7.55e-07 PS=3.24e-06
mXI20.XI3.MN_nand2 N_XI20.NET7_XI20.XI3.MN_nand2_d
+ N_XI20.NET6_XI20.XI3.MN_nand2_g N_XI20.XI3.NET6_XI20.XI3.MN_nand2_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=1.59e-12 AS=7.55e-13
+ PD=3.59e-06 PS=7.55e-07
mXI20.XI3.MM0 N_XI20.NET7_XI20.XI3.MM0_d N_CLK_BY_5_XI20.XI3.MM0_g
+ N_VDD_XI20.XI3.MM0_s N_VDD_XI272.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=7.55e-13
+ AS=1.22e-12 PD=7.55e-07 PS=3.22e-06
mXI20.XI3.MP_nand2 N_XI20.NET7_XI20.XI3.MP_nand2_d
+ N_XI20.NET6_XI20.XI3.MP_nand2_g N_VDD_XI20.XI3.MP_nand2_s N_VDD_XI272.MP_inv_b
+ P_18 L=1.8e-07 W=2e-06 AD=7.55e-13 AS=1.38e-12 PD=7.55e-07 PS=3.38e-06
mXI21.XI4.MM1 N_XI21.XI4.NET6_XI21.XI4.MM1_d N_CLK_BY_7_XI21.XI4.MM1_g
+ N_VSS_XI21.XI4.MM1_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=7.55e-13
+ AS=1.24e-12 PD=7.55e-07 PS=3.24e-06
mXI21.XI4.MN_nand2 N_XI21.NET7_XI21.XI4.MN_nand2_d
+ N_XI21.NET6_XI21.XI4.MN_nand2_g N_XI21.XI4.NET6_XI21.XI4.MN_nand2_s
+ N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=2e-06 AD=1.59e-12 AS=7.55e-13
+ PD=3.59e-06 PS=7.55e-07
mXI21.XI4.MM0 N_XI21.NET7_XI21.XI4.MM0_d N_CLK_BY_7_XI21.XI4.MM0_g
+ N_VDD_XI21.XI4.MM0_s N_VDD_XI252.MP_inv_b P_18 L=1.8e-07 W=2e-06 AD=7.55e-13
+ AS=1.22e-12 PD=7.55e-07 PS=3.22e-06
mXI21.XI4.MP_nand2 N_XI21.NET7_XI21.XI4.MP_nand2_d
+ N_XI21.NET6_XI21.XI4.MP_nand2_g N_VDD_XI21.XI4.MP_nand2_s N_VDD_XI252.MP_inv_b
+ P_18 L=1.8e-07 W=2e-06 AD=7.55e-13 AS=1.38e-12 PD=7.55e-07 PS=3.38e-06
mXI302.MN_inv N_CLK_BY_2_BAR2_XI302.MN_inv_d N_CLK_BY_2_XI302.MN_inv_g
+ N_VSS_XI302.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=4e-06 AD=3.2e-12
+ AS=3.3e-12 PD=5.6e-06 PS=5.65e-06
mXI302.MP_inv N_CLK_BY_2_BAR2_XI302.MP_inv_d N_CLK_BY_2_XI302.MP_inv_g
+ N_VDD_XI302.MP_inv_s N_VDD_XI302.MP_inv_b P_18 L=1.8e-07 W=1.2e-05 AD=9.72e-12
+ AS=1.068e-11 PD=1.362e-05 PS=1.378e-05
mXI312.MN_inv N_CLK_BY_1_BAR2_XI312.MN_inv_d N_CLK3_XI312.MN_inv_g
+ N_VSS_XI312.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=4e-06 AD=3.2e-12
+ AS=3.3e-12 PD=5.6e-06 PS=5.65e-06
mXI312.MP_inv N_CLK_BY_1_BAR2_XI312.MP_inv_d N_CLK3_XI312.MP_inv_g
+ N_VDD_XI312.MP_inv_s N_VDD_XI312.MP_inv_b P_18 L=1.8e-07 W=1.2e-05 AD=9.72e-12
+ AS=1.068e-11 PD=1.362e-05 PS=1.378e-05
mXI292.MN_inv N_CLK_BY_3_BAR2_XI292.MN_inv_d N_CLK_BY_3_XI292.MN_inv_g
+ N_VSS_XI292.MN_inv_s N_VSS_XI214.MN_inv_b N_18 L=1.8e-07 W=4e-06 AD=3.2e-12
+ AS=3.3e-12 PD=5.6e-06 PS=5.65e-06
mXI292.MP_inv N_CLK_BY_3_BAR2_XI292.MP_inv_d N_CLK_BY_3_XI292.MP_inv_g
+ N_VDD_XI292.MP_inv_s N_VDD_XI214.MP_inv_b P_18 L=1.8e-07 W=1.2e-05 AD=9.72e-12
+ AS=1.068e-11 PD=1.362e-05 PS=1.378e-05
*
.include "freqdiv4_2.pex.netlist.FREQDIV4.pxi"
*
.ends
*
*
